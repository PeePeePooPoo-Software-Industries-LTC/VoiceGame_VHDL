library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Empty for now, NIOS II Implementation branch.







-- More test



-- This line has no purpose, but I wanted to type it.