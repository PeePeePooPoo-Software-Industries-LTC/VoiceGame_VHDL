-- niosii_test_ci_inc_max_shorts.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosii_test_ci_inc_max_shorts is
	generic (
		SHARED_COMB_AND_MULTI : integer := 0
	);
	port (
		ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => '0'); --       ci_slave.dataa
		ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => '0'); --               .datab
		ci_slave_result           : out std_logic_vector(31 downto 0);                    --               .result
		comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- comb_ci_master.dataa
		comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    --               .datab
		comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => '0'); --               .result
		ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => '0');
		ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => '0');
		ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => '0');
		ci_slave_estatus          : in  std_logic                     := '0';
		ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => '0');
		ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => '0');
		ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => '0');
		ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => '0');
		ci_slave_multi_clk        : in  std_logic                     := '0';
		ci_slave_multi_clken      : in  std_logic                     := '0';
		ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => '0');
		ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => '0');
		ci_slave_multi_done       : out std_logic;
		ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => '0');
		ci_slave_multi_readra     : in  std_logic                     := '0';
		ci_slave_multi_readrb     : in  std_logic                     := '0';
		ci_slave_multi_reset      : in  std_logic                     := '0';
		ci_slave_multi_reset_req  : in  std_logic                     := '0';
		ci_slave_multi_result     : out std_logic_vector(31 downto 0);
		ci_slave_multi_start      : in  std_logic                     := '0';
		ci_slave_multi_writerc    : in  std_logic                     := '0';
		ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => '0');
		ci_slave_readra           : in  std_logic                     := '0';
		ci_slave_readrb           : in  std_logic                     := '0';
		ci_slave_writerc          : in  std_logic                     := '0';
		comb_ci_master_a          : out std_logic_vector(4 downto 0);
		comb_ci_master_b          : out std_logic_vector(4 downto 0);
		comb_ci_master_c          : out std_logic_vector(4 downto 0);
		comb_ci_master_estatus    : out std_logic;
		comb_ci_master_ipending   : out std_logic_vector(31 downto 0);
		comb_ci_master_n          : out std_logic_vector(7 downto 0);
		comb_ci_master_readra     : out std_logic;
		comb_ci_master_readrb     : out std_logic;
		comb_ci_master_writerc    : out std_logic;
		multi_ci_master_a         : out std_logic_vector(4 downto 0);
		multi_ci_master_b         : out std_logic_vector(4 downto 0);
		multi_ci_master_c         : out std_logic_vector(4 downto 0);
		multi_ci_master_clk       : out std_logic;
		multi_ci_master_clken     : out std_logic;
		multi_ci_master_dataa     : out std_logic_vector(31 downto 0);
		multi_ci_master_datab     : out std_logic_vector(31 downto 0);
		multi_ci_master_done      : in  std_logic                     := '0';
		multi_ci_master_n         : out std_logic_vector(7 downto 0);
		multi_ci_master_readra    : out std_logic;
		multi_ci_master_readrb    : out std_logic;
		multi_ci_master_reset     : out std_logic;
		multi_ci_master_reset_req : out std_logic;
		multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => '0');
		multi_ci_master_start     : out std_logic;
		multi_ci_master_writerc   : out std_logic
	);
end entity niosii_test_ci_inc_max_shorts;

architecture rtl of niosii_test_ci_inc_max_shorts is
	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_c
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0)                      -- c
		);
	end component altera_customins_master_translator;

begin

	shared_comb_and_multi_check : if SHARED_COMB_AND_MULTI /= 0 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	ci_inc_max_shorts : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 0
		)
		port map (
			ci_slave_dataa            => ci_slave_dataa,                     --       ci_slave.dataa
			ci_slave_datab            => ci_slave_datab,                     --               .datab
			ci_slave_result           => ci_slave_result,                    --               .result
			comb_ci_master_dataa      => comb_ci_master_dataa,               -- comb_ci_master.dataa
			comb_ci_master_datab      => comb_ci_master_datab,               --               .datab
			comb_ci_master_result     => comb_ci_master_result,              --               .result
			ci_slave_n                => "00000000",                         --    (terminated)
			ci_slave_readra           => '0',                                --    (terminated)
			ci_slave_readrb           => '0',                                --    (terminated)
			ci_slave_writerc          => '0',                                --    (terminated)
			ci_slave_a                => "00000",                            --    (terminated)
			ci_slave_b                => "00000",                            --    (terminated)
			ci_slave_c                => "00000",                            --    (terminated)
			ci_slave_ipending         => "00000000000000000000000000000000", --    (terminated)
			ci_slave_estatus          => '0',                                --    (terminated)
			ci_slave_multi_clk        => '0',                                --    (terminated)
			ci_slave_multi_reset      => '0',                                --    (terminated)
			ci_slave_multi_clken      => '0',                                --    (terminated)
			ci_slave_multi_reset_req  => '0',                                --    (terminated)
			ci_slave_multi_start      => '0',                                --    (terminated)
			ci_slave_multi_done       => open,                               --    (terminated)
			ci_slave_multi_dataa      => "00000000000000000000000000000000", --    (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000", --    (terminated)
			ci_slave_multi_result     => open,                               --    (terminated)
			ci_slave_multi_n          => "00000000",                         --    (terminated)
			ci_slave_multi_readra     => '0',                                --    (terminated)
			ci_slave_multi_readrb     => '0',                                --    (terminated)
			ci_slave_multi_writerc    => '0',                                --    (terminated)
			ci_slave_multi_a          => "00000",                            --    (terminated)
			ci_slave_multi_b          => "00000",                            --    (terminated)
			ci_slave_multi_c          => "00000",                            --    (terminated)
			comb_ci_master_n          => open,                               --    (terminated)
			comb_ci_master_readra     => open,                               --    (terminated)
			comb_ci_master_readrb     => open,                               --    (terminated)
			comb_ci_master_writerc    => open,                               --    (terminated)
			comb_ci_master_a          => open,                               --    (terminated)
			comb_ci_master_b          => open,                               --    (terminated)
			comb_ci_master_c          => open,                               --    (terminated)
			comb_ci_master_ipending   => open,                               --    (terminated)
			comb_ci_master_estatus    => open,                               --    (terminated)
			multi_ci_master_clk       => open,                               --    (terminated)
			multi_ci_master_reset     => open,                               --    (terminated)
			multi_ci_master_clken     => open,                               --    (terminated)
			multi_ci_master_reset_req => open,                               --    (terminated)
			multi_ci_master_start     => open,                               --    (terminated)
			multi_ci_master_done      => '0',                                --    (terminated)
			multi_ci_master_dataa     => open,                               --    (terminated)
			multi_ci_master_datab     => open,                               --    (terminated)
			multi_ci_master_result    => "00000000000000000000000000000000", --    (terminated)
			multi_ci_master_n         => open,                               --    (terminated)
			multi_ci_master_readra    => open,                               --    (terminated)
			multi_ci_master_readrb    => open,                               --    (terminated)
			multi_ci_master_writerc   => open,                               --    (terminated)
			multi_ci_master_a         => open,                               --    (terminated)
			multi_ci_master_b         => open,                               --    (terminated)
			multi_ci_master_c         => open                                --    (terminated)
		);

end architecture rtl; -- of niosii_test_ci_inc_max_shorts
