-- NIOSII_Test.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NIOSII_Test is
	port (
		audio_interface_ADCDAT                        : in    std_logic                     := '0';             --                        audio_interface.ADCDAT
		audio_interface_ADCLRCK                       : in    std_logic                     := '0';             --                                       .ADCLRCK
		audio_interface_BCLK                          : in    std_logic                     := '0';             --                                       .BCLK
		clk_clk                                       : in    std_logic                     := '0';             --                                    clk.clk
		pio_pixel_color_external_connection_export    : out   std_logic_vector(23 downto 0);                    --    pio_pixel_color_external_connection.export
		pio_pixel_position_external_connection_export : in    std_logic_vector(31 downto 0) := (others => '0'); -- pio_pixel_position_external_connection.export
		pio_request_external_connection_export        : in    std_logic                     := '0';             --        pio_request_external_connection.export
		reset_reset                                   : in    std_logic                     := '0';             --                                  reset.reset
		sdram_clk_clk                                 : out   std_logic;                                        --                              sdram_clk.clk
		sdram_wire_addr                               : out   std_logic_vector(11 downto 0);                    --                             sdram_wire.addr
		sdram_wire_ba                                 : out   std_logic;                                        --                                       .ba
		sdram_wire_cas_n                              : out   std_logic;                                        --                                       .cas_n
		sdram_wire_cke                                : out   std_logic;                                        --                                       .cke
		sdram_wire_cs_n                               : out   std_logic;                                        --                                       .cs_n
		sdram_wire_dq                                 : inout std_logic_vector(31 downto 0) := (others => '0'); --                                       .dq
		sdram_wire_dqm                                : out   std_logic_vector(3 downto 0);                     --                                       .dqm
		sdram_wire_ras_n                              : out   std_logic;                                        --                                       .ras_n
		sdram_wire_we_n                               : out   std_logic;                                        --                                       .we_n
		vga_CLK                                       : out   std_logic;                                        --                                    vga.CLK
		vga_HS                                        : out   std_logic;                                        --                                       .HS
		vga_VS                                        : out   std_logic;                                        --                                       .VS
		vga_BLANK                                     : out   std_logic;                                        --                                       .BLANK
		vga_SYNC                                      : out   std_logic;                                        --                                       .SYNC
		vga_R                                         : out   std_logic_vector(7 downto 0);                     --                                       .R
		vga_G                                         : out   std_logic_vector(7 downto 0);                     --                                       .G
		vga_B                                         : out   std_logic_vector(7 downto 0)                      --                                       .B
	);
end entity NIOSII_Test;

architecture rtl of NIOSII_Test is
	component NIOSII_Test_audio_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X'              -- export
		);
	end component NIOSII_Test_audio_0;

	component NIOSII_Test_audio_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component NIOSII_Test_audio_pll_0;

	component NIOSII_Test_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component NIOSII_Test_jtag_uart_0;

	component NIOSII_Test_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(20 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic;                                        -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component NIOSII_Test_new_sdram_controller_0;

	component NIOSII_Test_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(24 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component NIOSII_Test_nios2_gen2_0;

	component NIOSII_Test_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component NIOSII_Test_onchip_memory2_0;

	component NIOSII_Test_pio_pixel_color is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(23 downto 0)                     -- export
		);
	end component NIOSII_Test_pio_pixel_color;

	component NIOSII_Test_pio_pixel_position is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component NIOSII_Test_pio_pixel_position;

	component NIOSII_Test_pio_request is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOSII_Test_pio_request;

	component NIOSII_Test_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component NIOSII_Test_sys_sdram_pll_0;

	component NIOSII_Test_video_pixel_buffer_dma_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component NIOSII_Test_video_pixel_buffer_dma_0;

	component NIOSII_Test_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component NIOSII_Test_video_pll_0;

	component NIOSII_Test_video_vga_controller_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component NIOSII_Test_video_vga_controller_0;

	component NIOSII_Test_mm_interconnect_0 is
		port (
			audio_pll_0_audio_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			sys_sdram_pll_0_sys_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			video_pll_0_vga_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			audio_0_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			new_sdram_controller_0_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			onchip_memory2_0_reset1_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid                         : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                        : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_address       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest   : out std_logic;                                        -- waitrequest
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_read          : in  std_logic                     := 'X';             -- read
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid : out std_logic;                                        -- readdatavalid
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock          : in  std_logic                     := 'X';             -- lock
			audio_0_avalon_audio_slave_address                             : out std_logic_vector(1 downto 0);                     -- address
			audio_0_avalon_audio_slave_write                               : out std_logic;                                        -- write
			audio_0_avalon_audio_slave_read                                : out std_logic;                                        -- read
			audio_0_avalon_audio_slave_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_0_avalon_audio_slave_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			audio_0_avalon_audio_slave_chipselect                          : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                       : out std_logic;                                        -- chipselect
			new_sdram_controller_0_s1_address                              : out std_logic_vector(20 downto 0);                    -- address
			new_sdram_controller_0_s1_write                                : out std_logic;                                        -- write
			new_sdram_controller_0_s1_read                                 : out std_logic;                                        -- read
			new_sdram_controller_0_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			new_sdram_controller_0_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			new_sdram_controller_0_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			new_sdram_controller_0_s1_readdatavalid                        : in  std_logic                     := 'X';             -- readdatavalid
			new_sdram_controller_0_s1_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_chipselect                           : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                    : out std_logic_vector(16 downto 0);                    -- address
			onchip_memory2_0_s1_write                                      : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                      : out std_logic;                                        -- clken
			pio_pixel_color_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			pio_pixel_color_s1_write                                       : out std_logic;                                        -- write
			pio_pixel_color_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_pixel_color_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_pixel_color_s1_chipselect                                  : out std_logic;                                        -- chipselect
			pio_pixel_position_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			pio_pixel_position_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_request_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			pio_request_s1_write                                           : out std_logic;                                        -- write
			pio_request_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_request_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			pio_request_s1_chipselect                                      : out std_logic;                                        -- chipselect
			video_pixel_buffer_dma_0_avalon_control_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			video_pixel_buffer_dma_0_avalon_control_slave_write            : out std_logic;                                        -- write
			video_pixel_buffer_dma_0_avalon_control_slave_read             : out std_logic;                                        -- read
			video_pixel_buffer_dma_0_avalon_control_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_pixel_buffer_dma_0_avalon_control_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			video_pixel_buffer_dma_0_avalon_control_slave_byteenable       : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component NIOSII_Test_mm_interconnect_0;

	component NIOSII_Test_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component NIOSII_Test_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component niosii_test_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component niosii_test_rst_controller;

	component niosii_test_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component niosii_test_rst_controller_002;

	component niosii_test_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component niosii_test_rst_controller_003;

	signal video_pixel_buffer_dma_0_avalon_pixel_source_valid                         : std_logic;                     -- video_pixel_buffer_dma_0:stream_valid -> video_vga_controller_0:valid
	signal video_pixel_buffer_dma_0_avalon_pixel_source_data                          : std_logic_vector(29 downto 0); -- video_pixel_buffer_dma_0:stream_data -> video_vga_controller_0:data
	signal video_pixel_buffer_dma_0_avalon_pixel_source_ready                         : std_logic;                     -- video_vga_controller_0:ready -> video_pixel_buffer_dma_0:stream_ready
	signal video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket                 : std_logic;                     -- video_pixel_buffer_dma_0:stream_startofpacket -> video_vga_controller_0:startofpacket
	signal video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket                   : std_logic;                     -- video_pixel_buffer_dma_0:stream_endofpacket -> video_vga_controller_0:endofpacket
	signal audio_pll_0_audio_clk_clk                                                  : std_logic;                     -- audio_pll_0:audio_clk_clk -> [audio_0:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:audio_pll_0_audio_clk_clk, rst_controller:clk]
	signal sys_sdram_pll_0_sys_clk_clk                                                : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [audio_pll_0:ref_clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, pio_pixel_color:clk, pio_pixel_position:clk, pio_request:clk, rst_controller_001:clk, rst_controller_002:clk, rst_controller_003:clk, video_pll_0:ref_clk_clk]
	signal video_pll_0_vga_clk_clk                                                    : std_logic;                     -- video_pll_0:vga_clk_clk -> [mm_interconnect_0:video_pll_0_vga_clk_clk, rst_controller_004:clk, video_pixel_buffer_dma_0:clk, video_vga_controller_0:clk]
	signal video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest               : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma_0:master_waitrequest
	signal video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma_0:master_readdata
	signal video_pixel_buffer_dma_0_avalon_pixel_dma_master_address                   : std_logic_vector(31 downto 0); -- video_pixel_buffer_dma_0:master_address -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_address
	signal video_pixel_buffer_dma_0_avalon_pixel_dma_master_read                      : std_logic;                     -- video_pixel_buffer_dma_0:master_read -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_read
	signal video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid             : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma_0:master_readdatavalid
	signal video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock                      : std_logic;                     -- video_pixel_buffer_dma_0:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock
	signal nios2_gen2_0_data_master_readdata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                       : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                           : std_logic_vector(24 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                        : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                              : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                             : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                         : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                    : std_logic_vector(24 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                       : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_new_sdram_controller_0_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdata                       : std_logic_vector(31 downto 0); -- new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	signal mm_interconnect_0_new_sdram_controller_0_s1_waitrequest                    : std_logic;                     -- new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_new_sdram_controller_0_s1_address                        : std_logic_vector(20 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	signal mm_interconnect_0_new_sdram_controller_0_s1_read                           : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_read -> mm_interconnect_0_new_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> mm_interconnect_0_new_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid                  : std_logic;                     -- new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_new_sdram_controller_0_s1_write                          : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_write -> mm_interconnect_0_new_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                    : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                 : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                        : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                             : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                              : std_logic_vector(16 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_audio_0_avalon_audio_slave_chipselect                    : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_chipselect -> audio_0:chipselect
	signal mm_interconnect_0_audio_0_avalon_audio_slave_readdata                      : std_logic_vector(31 downto 0); -- audio_0:readdata -> mm_interconnect_0:audio_0_avalon_audio_slave_readdata
	signal mm_interconnect_0_audio_0_avalon_audio_slave_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_0_avalon_audio_slave_address -> audio_0:address
	signal mm_interconnect_0_audio_0_avalon_audio_slave_read                          : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_read -> audio_0:read
	signal mm_interconnect_0_audio_0_avalon_audio_slave_write                         : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_write -> audio_0:write
	signal mm_interconnect_0_audio_0_avalon_audio_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_0_avalon_audio_slave_writedata -> audio_0:writedata
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata   : std_logic_vector(31 downto 0); -- video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read       : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write      : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	signal mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                 : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                   : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                       : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_pio_pixel_position_s1_readdata                           : std_logic_vector(31 downto 0); -- pio_pixel_position:readdata -> mm_interconnect_0:pio_pixel_position_s1_readdata
	signal mm_interconnect_0_pio_pixel_position_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_pixel_position_s1_address -> pio_pixel_position:address
	signal mm_interconnect_0_pio_request_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:pio_request_s1_chipselect -> pio_request:chipselect
	signal mm_interconnect_0_pio_request_s1_readdata                                  : std_logic_vector(31 downto 0); -- pio_request:readdata -> mm_interconnect_0:pio_request_s1_readdata
	signal mm_interconnect_0_pio_request_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_request_s1_address -> pio_request:address
	signal mm_interconnect_0_pio_request_s1_write                                     : std_logic;                     -- mm_interconnect_0:pio_request_s1_write -> mm_interconnect_0_pio_request_s1_write:in
	signal mm_interconnect_0_pio_request_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_request_s1_writedata -> pio_request:writedata
	signal mm_interconnect_0_pio_pixel_color_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:pio_pixel_color_s1_chipselect -> pio_pixel_color:chipselect
	signal mm_interconnect_0_pio_pixel_color_s1_readdata                              : std_logic_vector(31 downto 0); -- pio_pixel_color:readdata -> mm_interconnect_0:pio_pixel_color_s1_readdata
	signal mm_interconnect_0_pio_pixel_color_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_pixel_color_s1_address -> pio_pixel_color:address
	signal mm_interconnect_0_pio_pixel_color_s1_write                                 : std_logic;                     -- mm_interconnect_0:pio_pixel_color_s1_write -> mm_interconnect_0_pio_pixel_color_s1_write:in
	signal mm_interconnect_0_pio_pixel_color_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_pixel_color_s1_writedata -> pio_pixel_color:writedata
	signal irq_mapper_receiver1_irq                                                   : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                   : std_logic;                     -- pio_request:irq -> irq_mapper:receiver2_irq
	signal nios2_gen2_0_irq_irq                                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver0_irq                                                   : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                              : std_logic_vector(0 downto 0);  -- audio_0:irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                             : std_logic;                     -- rst_controller:reset_out -> [audio_0:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:audio_0_reset_reset_bridge_in_reset_reset]
	signal audio_pll_0_reset_source_reset                                             : std_logic;                     -- audio_pll_0:reset_source_reset -> rst_controller:reset_in0
	signal rst_controller_001_reset_out_reset                                         : std_logic;                     -- rst_controller_001:reset_out -> [audio_pll_0:ref_reset_reset, mm_interconnect_0:new_sdram_controller_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, video_pll_0:ref_reset_reset]
	signal sys_sdram_pll_0_reset_source_reset                                         : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> [rst_controller_001:reset_in0, rst_controller_003:reset_in1]
	signal rst_controller_002_reset_out_reset                                         : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_002_reset_out_reset_req                                     : std_logic;                     -- rst_controller_002:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                                     : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal rst_controller_003_reset_out_reset                                         : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	signal rst_controller_003_reset_out_reset_req                                     : std_logic;                     -- rst_controller_003:reset_req -> onchip_memory2_0:reset_req
	signal rst_controller_004_reset_out_reset                                         : std_logic;                     -- rst_controller_004:reset_out -> [mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, video_pixel_buffer_dma_0:reset, video_vga_controller_0:reset]
	signal video_pll_0_reset_source_reset                                             : std_logic;                     -- video_pll_0:reset_source_reset -> rst_controller_004:reset_in0
	signal mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv                 : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_read:inv -> new_sdram_controller_0:az_rd_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv           : std_logic_vector(3 downto 0);  -- mm_interconnect_0_new_sdram_controller_0_s1_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_write:inv -> new_sdram_controller_0:az_wr_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv             : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv            : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_pio_request_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_pio_request_s1_write:inv -> pio_request:write_n
	signal mm_interconnect_0_pio_pixel_color_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_pio_pixel_color_s1_write:inv -> pio_pixel_color:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [new_sdram_controller_0:reset_n, pio_pixel_color:reset_n, pio_pixel_position:reset_n, pio_request:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [jtag_uart_0:rst_n, nios2_gen2_0:reset_n]

begin

	audio_0 : component NIOSII_Test_audio_0
		port map (
			clk         => audio_pll_0_audio_clk_clk,                               --                clk.clk
			reset       => rst_controller_reset_out_reset,                          --              reset.reset
			address     => mm_interconnect_0_audio_0_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_0_audio_0_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_0_audio_0_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,   --                   .readdata
			irq         => irq_synchronizer_receiver_irq(0),                        --          interrupt.irq
			AUD_ADCDAT  => audio_interface_ADCDAT,                                  -- external_interface.export
			AUD_ADCLRCK => audio_interface_ADCLRCK,                                 --                   .export
			AUD_BCLK    => audio_interface_BCLK                                     --                   .export
		);

	audio_pll_0 : component NIOSII_Test_audio_pll_0
		port map (
			ref_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			audio_clk_clk      => audio_pll_0_audio_clk_clk,          --    audio_clk.clk
			reset_source_reset => audio_pll_0_reset_source_reset      -- reset_source.reset
		);

	jtag_uart_0 : component NIOSII_Test_jtag_uart_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                     --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	new_sdram_controller_0 : component NIOSII_Test_new_sdram_controller_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => mm_interconnect_0_new_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_new_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_new_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                                  --  wire.export
			zs_ba          => sdram_wire_ba,                                                    --      .export
			zs_cas_n       => sdram_wire_cas_n,                                                 --      .export
			zs_cke         => sdram_wire_cke,                                                   --      .export
			zs_cs_n        => sdram_wire_cs_n,                                                  --      .export
			zs_dq          => sdram_wire_dq,                                                    --      .export
			zs_dqm         => sdram_wire_dqm,                                                   --      .export
			zs_ras_n       => sdram_wire_ras_n,                                                 --      .export
			zs_we_n        => sdram_wire_we_n                                                   --      .export
		);

	nios2_gen2_0 : component NIOSII_Test_nios2_gen2_0
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                                --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component NIOSII_Test_onchip_memory2_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                      --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_003_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_003_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	pio_pixel_color : component NIOSII_Test_pio_pixel_color
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_pio_pixel_color_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_pixel_color_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_pixel_color_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_pixel_color_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_pixel_color_s1_readdata,        --                    .readdata
			out_port   => pio_pixel_color_external_connection_export            -- external_connection.export
		);

	pio_pixel_position : component NIOSII_Test_pio_pixel_position
		port map (
			clk      => sys_sdram_pll_0_sys_clk_clk,                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,     --               reset.reset_n
			address  => mm_interconnect_0_pio_pixel_position_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_pixel_position_s1_readdata, --                    .readdata
			in_port  => pio_pixel_position_external_connection_export     -- external_connection.export
		);

	pio_request : component NIOSII_Test_pio_request
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_request_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_request_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_request_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_request_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_request_s1_readdata,        --                    .readdata
			in_port    => pio_request_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                          --                 irq.irq
		);

	sys_sdram_pll_0 : component NIOSII_Test_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => reset_reset,                        --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	video_pixel_buffer_dma_0 : component NIOSII_Test_video_pixel_buffer_dma_0
		port map (
			clk                  => video_pll_0_vga_clk_clk,                                                    --                     clk.clk
			reset                => rst_controller_004_reset_out_reset,                                         --                   reset.reset
			master_readdatavalid => video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid,             -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest,               --                        .waitrequest
			master_address       => video_pixel_buffer_dma_0_avalon_pixel_dma_master_address,                   --                        .address
			master_arbiterlock   => video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock,                      --                        .lock
			master_read          => video_pixel_buffer_dma_0_avalon_pixel_dma_master_read,                      --                        .read
			master_readdata      => video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata,                  --                        .readdata
			slave_address        => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address,    --    avalon_control_slave.address
			slave_byteenable     => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable, --                        .byteenable
			slave_read           => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read,       --                        .read
			slave_write          => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write,      --                        .write
			slave_writedata      => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata,  --                        .writedata
			slave_readdata       => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata,   --                        .readdata
			stream_ready         => video_pixel_buffer_dma_0_avalon_pixel_source_ready,                         --     avalon_pixel_source.ready
			stream_startofpacket => video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket,                 --                        .startofpacket
			stream_endofpacket   => video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket,                   --                        .endofpacket
			stream_valid         => video_pixel_buffer_dma_0_avalon_pixel_source_valid,                         --                        .valid
			stream_data          => video_pixel_buffer_dma_0_avalon_pixel_source_data                           --                        .data
		);

	video_pll_0 : component NIOSII_Test_video_pll_0
		port map (
			ref_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			vga_clk_clk        => video_pll_0_vga_clk_clk,            --      vga_clk.clk
			reset_source_reset => video_pll_0_reset_source_reset      -- reset_source.reset
		);

	video_vga_controller_0 : component NIOSII_Test_video_vga_controller_0
		port map (
			clk           => video_pll_0_vga_clk_clk,                                    --                clk.clk
			reset         => rst_controller_004_reset_out_reset,                         --              reset.reset
			data          => video_pixel_buffer_dma_0_avalon_pixel_source_data,          --    avalon_vga_sink.data
			startofpacket => video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket, --                   .startofpacket
			endofpacket   => video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket,   --                   .endofpacket
			valid         => video_pixel_buffer_dma_0_avalon_pixel_source_valid,         --                   .valid
			ready         => video_pixel_buffer_dma_0_avalon_pixel_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                                    -- external_interface.export
			VGA_HS        => vga_HS,                                                     --                   .export
			VGA_VS        => vga_VS,                                                     --                   .export
			VGA_BLANK     => vga_BLANK,                                                  --                   .export
			VGA_SYNC      => vga_SYNC,                                                   --                   .export
			VGA_R         => vga_R,                                                      --                   .export
			VGA_G         => vga_G,                                                      --                   .export
			VGA_B         => vga_B                                                       --                   .export
		);

	mm_interconnect_0 : component NIOSII_Test_mm_interconnect_0
		port map (
			audio_pll_0_audio_clk_clk                                      => audio_pll_0_audio_clk_clk,                                                  --                                audio_pll_0_audio_clk.clk
			sys_sdram_pll_0_sys_clk_clk                                    => sys_sdram_pll_0_sys_clk_clk,                                                --                              sys_sdram_pll_0_sys_clk.clk
			video_pll_0_vga_clk_clk                                        => video_pll_0_vga_clk_clk,                                                    --                                  video_pll_0_vga_clk.clk
			audio_0_reset_reset_bridge_in_reset_reset                      => rst_controller_reset_out_reset,                                             --                  audio_0_reset_reset_bridge_in_reset.reset
			new_sdram_controller_0_reset_reset_bridge_in_reset_reset       => rst_controller_001_reset_out_reset,                                         --   new_sdram_controller_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                 => rst_controller_002_reset_out_reset,                                         --             nios2_gen2_0_reset_reset_bridge_in_reset.reset
			onchip_memory2_0_reset1_reset_bridge_in_reset_reset            => rst_controller_003_reset_out_reset,                                         --        onchip_memory2_0_reset1_reset_bridge_in_reset.reset
			video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset     => rst_controller_004_reset_out_reset,                                         -- video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                               => nios2_gen2_0_data_master_address,                                           --                             nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                           => nios2_gen2_0_data_master_waitrequest,                                       --                                                     .waitrequest
			nios2_gen2_0_data_master_byteenable                            => nios2_gen2_0_data_master_byteenable,                                        --                                                     .byteenable
			nios2_gen2_0_data_master_read                                  => nios2_gen2_0_data_master_read,                                              --                                                     .read
			nios2_gen2_0_data_master_readdata                              => nios2_gen2_0_data_master_readdata,                                          --                                                     .readdata
			nios2_gen2_0_data_master_readdatavalid                         => nios2_gen2_0_data_master_readdatavalid,                                     --                                                     .readdatavalid
			nios2_gen2_0_data_master_write                                 => nios2_gen2_0_data_master_write,                                             --                                                     .write
			nios2_gen2_0_data_master_writedata                             => nios2_gen2_0_data_master_writedata,                                         --                                                     .writedata
			nios2_gen2_0_data_master_debugaccess                           => nios2_gen2_0_data_master_debugaccess,                                       --                                                     .debugaccess
			nios2_gen2_0_instruction_master_address                        => nios2_gen2_0_instruction_master_address,                                    --                      nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                    => nios2_gen2_0_instruction_master_waitrequest,                                --                                                     .waitrequest
			nios2_gen2_0_instruction_master_read                           => nios2_gen2_0_instruction_master_read,                                       --                                                     .read
			nios2_gen2_0_instruction_master_readdata                       => nios2_gen2_0_instruction_master_readdata,                                   --                                                     .readdata
			nios2_gen2_0_instruction_master_readdatavalid                  => nios2_gen2_0_instruction_master_readdatavalid,                              --                                                     .readdatavalid
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_address       => video_pixel_buffer_dma_0_avalon_pixel_dma_master_address,                   --     video_pixel_buffer_dma_0_avalon_pixel_dma_master.address
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest   => video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest,               --                                                     .waitrequest
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_read          => video_pixel_buffer_dma_0_avalon_pixel_dma_master_read,                      --                                                     .read
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata      => video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata,                  --                                                     .readdata
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid => video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid,             --                                                     .readdatavalid
			video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock          => video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock,                      --                                                     .lock
			audio_0_avalon_audio_slave_address                             => mm_interconnect_0_audio_0_avalon_audio_slave_address,                       --                           audio_0_avalon_audio_slave.address
			audio_0_avalon_audio_slave_write                               => mm_interconnect_0_audio_0_avalon_audio_slave_write,                         --                                                     .write
			audio_0_avalon_audio_slave_read                                => mm_interconnect_0_audio_0_avalon_audio_slave_read,                          --                                                     .read
			audio_0_avalon_audio_slave_readdata                            => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,                      --                                                     .readdata
			audio_0_avalon_audio_slave_writedata                           => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,                     --                                                     .writedata
			audio_0_avalon_audio_slave_chipselect                          => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect,                    --                                                     .chipselect
			jtag_uart_0_avalon_jtag_slave_address                          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                    --                        jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                      --                                                     .write
			jtag_uart_0_avalon_jtag_slave_read                             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                       --                                                     .read
			jtag_uart_0_avalon_jtag_slave_readdata                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                   --                                                     .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,                  --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,                --                                                     .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,                 --                                                     .chipselect
			new_sdram_controller_0_s1_address                              => mm_interconnect_0_new_sdram_controller_0_s1_address,                        --                            new_sdram_controller_0_s1.address
			new_sdram_controller_0_s1_write                                => mm_interconnect_0_new_sdram_controller_0_s1_write,                          --                                                     .write
			new_sdram_controller_0_s1_read                                 => mm_interconnect_0_new_sdram_controller_0_s1_read,                           --                                                     .read
			new_sdram_controller_0_s1_readdata                             => mm_interconnect_0_new_sdram_controller_0_s1_readdata,                       --                                                     .readdata
			new_sdram_controller_0_s1_writedata                            => mm_interconnect_0_new_sdram_controller_0_s1_writedata,                      --                                                     .writedata
			new_sdram_controller_0_s1_byteenable                           => mm_interconnect_0_new_sdram_controller_0_s1_byteenable,                     --                                                     .byteenable
			new_sdram_controller_0_s1_readdatavalid                        => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,                  --                                                     .readdatavalid
			new_sdram_controller_0_s1_waitrequest                          => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,                    --                                                     .waitrequest
			new_sdram_controller_0_s1_chipselect                           => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,                     --                                                     .chipselect
			nios2_gen2_0_debug_mem_slave_address                           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                     --                         nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                       --                                                     .write
			nios2_gen2_0_debug_mem_slave_read                              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                        --                                                     .read
			nios2_gen2_0_debug_mem_slave_readdata                          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                    --                                                     .readdata
			nios2_gen2_0_debug_mem_slave_writedata                         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,                   --                                                     .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,                  --                                                     .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,                 --                                                     .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,                 --                                                     .debugaccess
			onchip_memory2_0_s1_address                                    => mm_interconnect_0_onchip_memory2_0_s1_address,                              --                                  onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                      => mm_interconnect_0_onchip_memory2_0_s1_write,                                --                                                     .write
			onchip_memory2_0_s1_readdata                                   => mm_interconnect_0_onchip_memory2_0_s1_readdata,                             --                                                     .readdata
			onchip_memory2_0_s1_writedata                                  => mm_interconnect_0_onchip_memory2_0_s1_writedata,                            --                                                     .writedata
			onchip_memory2_0_s1_byteenable                                 => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                           --                                                     .byteenable
			onchip_memory2_0_s1_chipselect                                 => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                           --                                                     .chipselect
			onchip_memory2_0_s1_clken                                      => mm_interconnect_0_onchip_memory2_0_s1_clken,                                --                                                     .clken
			pio_pixel_color_s1_address                                     => mm_interconnect_0_pio_pixel_color_s1_address,                               --                                   pio_pixel_color_s1.address
			pio_pixel_color_s1_write                                       => mm_interconnect_0_pio_pixel_color_s1_write,                                 --                                                     .write
			pio_pixel_color_s1_readdata                                    => mm_interconnect_0_pio_pixel_color_s1_readdata,                              --                                                     .readdata
			pio_pixel_color_s1_writedata                                   => mm_interconnect_0_pio_pixel_color_s1_writedata,                             --                                                     .writedata
			pio_pixel_color_s1_chipselect                                  => mm_interconnect_0_pio_pixel_color_s1_chipselect,                            --                                                     .chipselect
			pio_pixel_position_s1_address                                  => mm_interconnect_0_pio_pixel_position_s1_address,                            --                                pio_pixel_position_s1.address
			pio_pixel_position_s1_readdata                                 => mm_interconnect_0_pio_pixel_position_s1_readdata,                           --                                                     .readdata
			pio_request_s1_address                                         => mm_interconnect_0_pio_request_s1_address,                                   --                                       pio_request_s1.address
			pio_request_s1_write                                           => mm_interconnect_0_pio_request_s1_write,                                     --                                                     .write
			pio_request_s1_readdata                                        => mm_interconnect_0_pio_request_s1_readdata,                                  --                                                     .readdata
			pio_request_s1_writedata                                       => mm_interconnect_0_pio_request_s1_writedata,                                 --                                                     .writedata
			pio_request_s1_chipselect                                      => mm_interconnect_0_pio_request_s1_chipselect,                                --                                                     .chipselect
			video_pixel_buffer_dma_0_avalon_control_slave_address          => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address,    --        video_pixel_buffer_dma_0_avalon_control_slave.address
			video_pixel_buffer_dma_0_avalon_control_slave_write            => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write,      --                                                     .write
			video_pixel_buffer_dma_0_avalon_control_slave_read             => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read,       --                                                     .read
			video_pixel_buffer_dma_0_avalon_control_slave_readdata         => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata,   --                                                     .readdata
			video_pixel_buffer_dma_0_avalon_control_slave_writedata        => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata,  --                                                     .writedata
			video_pixel_buffer_dma_0_avalon_control_slave_byteenable       => mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable  --                                                     .byteenable
		);

	irq_mapper : component NIOSII_Test_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => audio_pll_0_audio_clk_clk,          --       receiver_clk.clk
			sender_clk     => sys_sdram_pll_0_sys_clk_clk,        --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	rst_controller : component niosii_test_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => audio_pll_0_reset_source_reset, -- reset_in0.reset
			clk            => audio_pll_0_audio_clk_clk,      --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component niosii_test_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_0_reset_source_reset, -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component niosii_test_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component niosii_test_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => sys_sdram_pll_0_reset_source_reset,     -- reset_in1.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_003_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_004 : component niosii_test_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => video_pll_0_reset_source_reset,     -- reset_in0.reset
			clk            => video_pll_0_vga_clk_clk,            --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_read;

	mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_write;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_pio_request_s1_write_ports_inv <= not mm_interconnect_0_pio_request_s1_write;

	mm_interconnect_0_pio_pixel_color_s1_write_ports_inv <= not mm_interconnect_0_pio_pixel_color_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of NIOSII_Test
